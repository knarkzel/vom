module character

// Based on https://docs.rs/nom/7.1.0/nom/character/index.html

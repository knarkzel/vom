module vom

fn test_alpha0() {
	// parser := is_a('123456789ABCDEF')
	// rest, output := parser('DEADBEEF and others') ?
	// assert output == 'DEADBEEF'
	// assert rest == ' and others'
}

module vom

// Based on https://docs.rs/nom/7.1.3/nom/number/complete/index.html

module vom

fn test_dummy() ? {
	assert 1 + 1 == 2
}

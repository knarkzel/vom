module vom

// Based on https://docs.rs/nom/7.1.0/nom/combinator/index.html

module vom

fn test_method() ? {
    assert 1 + 1 == 2
}

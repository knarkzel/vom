module vom

fn branch_test() ? {
}

fn permutation_test() ? {
}
